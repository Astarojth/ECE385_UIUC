// It's a full adder, which can also generate the p (propagating logic) and g (generating logic).


