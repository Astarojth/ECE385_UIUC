// It's a 4-bit carry lookahead adder.

